module AON_BUF_X1(A, Z);
  input A;
  output Z;
endmodule

module AON_BUF_X2(A, Z);
  input A;
  output Z;
endmodule

module AON_BUF_X4(A, Z);
  input A;
  output Z;
endmodule

module AON_INV_X1(A, Z);
  input A;
  output Z;
endmodule

module AON_INV_X2(A, Z);
  input A;
  output Z;
endmodule

module AON_INV_X4(A, Z);
  input A;
  output Z;
endmodule

module HEADER_OE_X1(SLEEP, SLEEPOUT);
  input SLEEP;
  output SLEEPOUT;
endmodule

module HEADER_OE_X2(SLEEP, SLEEPOUT);
  input SLEEP;
  output SLEEPOUT;
endmodule

module HEADER_OE_X4(SLEEP, SLEEPOUT);
  input SLEEP;
  output SLEEPOUT;
endmodule

module HEADER_X1(SLEEP);
  input SLEEP;
endmodule

module HEADER_X2(SLEEP);
  input SLEEP;
endmodule

module HEADER_X4(SLEEP);
  input SLEEP;
endmodule

module ISO_FENCE0N_X1(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE0N_X2(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE0N_X4(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE0_X1(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE0_X2(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE0_X4(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1N_X1(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1N_X2(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1N_X4(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1_X1(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1_X2(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module ISO_FENCE1_X4(A, EN, Z);
  input A;
  input EN;
  output Z;
endmodule

module LS_HLEN_X1(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_HLEN_X2(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_HLEN_X4(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_HL_X1(A, Z);
  input A;
  output Z;
endmodule

module LS_HL_X2(A, Z);
  input A;
  output Z;
endmodule

module LS_HL_X4(A, Z);
  input A;
  output Z;
endmodule

module LS_LHEN_X1(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_LHEN_X2(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_LHEN_X4(A, ISOLN, Z);
  input A;
  input ISOLN;
  output Z;
endmodule

module LS_LH_X1(A, Z);
  input A;
  output Z;
endmodule

module LS_LH_X2(A, Z);
  input A;
  output Z;
endmodule

module LS_LH_X4(A, Z);
  input A;
  output Z;
endmodule
